module dut_top (
   input CLK,
   input RST
);
   top DUT(.*);
   mult_top MULT_DUT(.*);

endmodule//dut_top
