// program test;
//    class regfile_random_item;
//       rand logic [ 31 : 0 ] data1;
//       rand logic [ 31 : 0 ] data2;
//       rand logic [ 4 : 0 ] addr1;
//       rand logic [ 4 : 0 ] addr2;
//    
//       function new();
//       endfunction
//    
//    endclass
//    
//    class regfile_random;
//       regfile_random_item rrr = new();
//    
//       function body();
//          rrr.randomize();
//       endfunction
//    
//    endclass
// endprogram
class a;
endclass
