parameter DATA_WIDTH=32;
parameter REG_ADDR_WIDTH=5;
