module dut_top (
   input CLK,
   input RST
);
   top DUT(.*);

endmodule//dut_top
